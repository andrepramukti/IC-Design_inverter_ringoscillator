magic
tech sky130A
magscale 1 2
timestamp 1729221103
<< nwell >>
rect -303 -898 951 2173
<< nsubdiff >>
rect -140 2003 -80 2037
rect 730 2003 786 2037
rect -140 1977 -106 2003
rect 752 1977 786 2003
rect -140 -742 -106 -716
rect 752 -742 786 -716
rect -140 -776 -80 -742
rect 730 -776 786 -742
<< nsubdiffcont >>
rect -80 2003 730 2037
rect -140 -716 -106 1977
rect 752 -716 786 1977
rect -80 -776 730 -742
<< poly >>
rect -59 1961 36 1977
rect -59 1927 -43 1961
rect -9 1927 36 1961
rect -59 1911 36 1927
rect 6 1876 36 1911
rect 610 1965 705 1981
rect 610 1931 655 1965
rect 689 1931 705 1965
rect 610 1915 705 1931
rect 610 1906 640 1915
rect 94 1283 294 1383
rect -59 1267 36 1283
rect -59 1233 -43 1267
rect -9 1233 36 1267
rect -59 1217 36 1233
rect 6 1182 36 1217
rect 610 1271 705 1287
rect 610 1237 655 1271
rect 689 1237 705 1271
rect 610 1221 705 1237
rect 610 1186 640 1221
rect 94 588 552 690
rect 6 61 36 96
rect -59 45 36 61
rect -59 11 -43 45
rect -9 11 36 45
rect -59 -5 36 11
rect 610 58 640 93
rect 610 42 705 58
rect 610 8 655 42
rect 689 8 705 42
rect 352 -106 552 -4
rect 610 -8 705 8
rect 5 -654 36 -628
rect -59 -670 36 -654
rect -59 -704 -43 -670
rect -9 -704 36 -670
rect -59 -720 36 -704
rect 610 -645 640 -610
rect 610 -661 705 -645
rect 610 -695 655 -661
rect 689 -695 705 -661
rect 610 -711 705 -695
<< polycont >>
rect -43 1927 -9 1961
rect 655 1931 689 1965
rect -43 1233 -9 1267
rect 655 1237 689 1271
rect -43 11 -9 45
rect 655 8 689 42
rect -43 -704 -9 -670
rect 655 -695 689 -661
<< locali >>
rect -140 2003 -80 2037
rect 730 2003 786 2037
rect -140 1977 -106 2003
rect 752 1977 786 2003
rect -59 1927 -43 1961
rect -9 1927 7 1961
rect 639 1931 655 1965
rect 689 1931 705 1965
rect -40 1876 -6 1927
rect 652 1879 686 1931
rect -38 1872 -8 1876
rect 656 1870 686 1879
rect -59 1233 -43 1267
rect -9 1233 7 1267
rect 639 1237 655 1271
rect 689 1237 705 1271
rect -40 1182 -6 1233
rect 652 1186 686 1237
rect -38 1178 -6 1182
rect 654 1176 686 1186
rect -40 45 -6 100
rect 656 93 686 102
rect -59 11 -43 45
rect -9 11 7 45
rect 652 42 686 93
rect 639 8 655 42
rect 689 8 705 42
rect 652 -205 686 -154
rect -38 -606 -6 -590
rect -40 -670 -6 -606
rect 652 -661 686 -590
rect -59 -704 -43 -670
rect -9 -704 7 -670
rect 639 -695 655 -661
rect 689 -695 705 -661
rect -140 -742 -106 -716
rect 752 -742 786 -716
rect -140 -776 -80 -742
rect 730 -776 786 -742
<< viali >>
rect 655 2003 689 2037
rect -43 1927 -9 1961
rect 655 1931 689 1965
rect 306 1492 340 1868
rect -43 1233 -9 1267
rect 655 1237 689 1271
rect 306 798 340 1174
rect 306 104 340 480
rect -43 11 -9 45
rect 655 8 689 42
rect 306 -590 340 -214
rect -43 -704 -9 -670
rect 655 -695 689 -661
rect -43 -776 -9 -742
<< metal1 >>
rect 643 2037 701 2043
rect 643 2003 655 2037
rect 689 2003 701 2037
rect -55 1961 3 1967
rect -55 1927 -43 1961
rect -9 1927 3 1961
rect -55 1921 3 1927
rect 643 1965 701 2003
rect 643 1931 655 1965
rect 689 1931 701 1965
rect 643 1925 701 1931
rect -44 1870 -4 1921
rect -60 1490 -50 1870
rect 2 1868 12 1870
rect 300 1868 346 1880
rect 650 1874 690 1925
rect 2 1492 82 1868
rect 300 1492 306 1868
rect 340 1492 346 1868
rect 564 1492 686 1868
rect 2 1490 12 1492
rect 300 1438 346 1492
rect 561 1438 599 1492
rect 300 1400 599 1438
rect 300 1393 559 1400
rect -55 1267 3 1273
rect -55 1233 -43 1267
rect -9 1233 3 1267
rect -55 1227 3 1233
rect -44 1182 3 1227
rect -40 1174 3 1182
rect 300 1174 346 1393
rect 643 1271 701 1277
rect 643 1237 655 1271
rect 689 1237 701 1271
rect 643 1231 701 1237
rect 650 1186 690 1231
rect -40 798 38 1174
rect 90 798 100 1174
rect 300 798 306 1174
rect 340 798 346 1174
rect 53 556 144 574
rect 48 540 144 556
rect 48 492 82 540
rect -48 102 98 492
rect 300 480 346 798
rect 554 788 688 1182
rect 564 740 598 788
rect 512 704 598 740
rect 300 104 306 480
rect 340 104 346 480
rect 546 104 556 480
rect 608 104 686 480
rect -44 51 -4 96
rect -55 45 3 51
rect -55 11 -43 45
rect -9 11 3 45
rect -55 5 3 11
rect 300 -117 346 104
rect 650 48 690 93
rect 643 42 701 48
rect 643 8 655 42
rect 689 8 701 42
rect 643 2 701 8
rect 42 -162 346 -117
rect 628 -154 688 -92
rect 42 -214 87 -162
rect 300 -214 346 -162
rect 643 -207 689 -154
rect 637 -214 647 -207
rect -4 -590 82 -214
rect 300 -590 306 -214
rect 340 -590 346 -214
rect 564 -269 647 -214
rect 716 -269 726 -207
rect 564 -590 650 -269
rect 706 -590 716 -269
rect 300 -602 346 -590
rect 650 -594 688 -593
rect -41 -641 -5 -602
rect -44 -664 -4 -641
rect 650 -655 690 -594
rect 643 -661 701 -655
rect -55 -670 3 -664
rect -55 -704 -43 -670
rect -9 -704 3 -670
rect 643 -695 655 -661
rect 689 -695 701 -661
rect 643 -701 701 -695
rect -55 -742 3 -704
rect -55 -776 -43 -742
rect -9 -776 3 -742
rect -55 -782 3 -776
<< via1 >>
rect -50 1490 2 1870
rect 38 798 90 1174
rect 556 104 608 480
rect 647 -269 716 -207
rect 650 -590 706 -269
<< metal2 >>
rect -50 1870 2 1880
rect -50 1480 2 1490
rect -44 1373 -4 1480
rect -44 1364 14 1373
rect -44 1308 -42 1364
rect -44 1299 14 1308
rect 628 1366 710 1382
rect 628 1306 638 1366
rect 698 1306 710 1366
rect -44 -21 -4 1299
rect 628 1290 710 1306
rect 38 1174 90 1184
rect 90 798 92 800
rect 38 788 92 798
rect 40 669 92 788
rect 552 669 606 670
rect 40 617 606 669
rect 552 490 606 617
rect 552 480 608 490
rect 556 94 608 104
rect -54 -30 6 -21
rect 650 -23 686 1290
rect 630 -30 686 -23
rect -54 -99 6 -90
rect 628 -32 688 -30
rect 628 -88 630 -32
rect 686 -88 688 -32
rect 628 -197 688 -88
rect 628 -206 716 -197
rect 647 -207 716 -206
rect 647 -279 650 -269
rect 706 -279 716 -269
rect 650 -600 706 -590
<< via2 >>
rect -42 1308 14 1364
rect 638 1306 698 1366
rect -54 -90 6 -30
rect 630 -88 686 -32
<< metal3 >>
rect -47 1366 19 1369
rect 633 1366 703 1371
rect -47 1364 638 1366
rect -47 1308 -42 1364
rect 14 1308 638 1364
rect -47 1306 638 1308
rect 698 1306 703 1366
rect -47 1303 19 1306
rect 633 1301 703 1306
rect -59 -30 11 -25
rect 625 -30 691 -27
rect -59 -90 -54 -30
rect 6 -32 691 -30
rect 6 -88 630 -32
rect 686 -88 691 -32
rect 6 -90 691 -88
rect -59 -95 11 -90
rect 625 -93 691 -90
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729147922
transform 1 0 625 0 1 1680
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729147922
transform 1 0 21 0 1 292
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729147922
transform 1 0 625 0 1 986
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729147922
transform 1 0 21 0 1 986
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729147922
transform 1 0 21 0 1 1680
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729147922
transform 1 0 625 0 1 292
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_8
timestamp 1729147922
transform 1 0 21 0 1 -402
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_9
timestamp 1729147922
transform 1 0 625 0 1 -402
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729147922
transform 1 0 323 0 1 1680
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729147922
transform 1 0 323 0 1 986
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729147922
transform 1 0 323 0 1 292
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729147922
transform 1 0 323 0 1 -402
box -323 -300 323 300
<< labels >>
flabel metal1 668 1994 668 1994 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal2 664 622 664 622 0 FreeSans 160 0 0 0 D5
port 1 nsew
flabel metal1 584 746 584 746 0 FreeSans 160 0 0 0 D2
port 2 nsew
flabel metal2 64 640 64 640 0 FreeSans 160 0 0 0 D1
port 3 nsew
<< end >>
